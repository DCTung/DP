module IDEXBuffer()
